/*
:name: integer_signed_bit
:description: bit signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
bit signed v;
endmodule