/*
:name: bufif1
:description: The 'bufif1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit bufif1;
endmodule