/*
:name: first_match
:description: The 'first_match' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit first_match;
endmodule