/*
:name: net_wand
:description: wand net test
:should_fail: 0
:tags: 6.6.3
*/
module top();
wand v;
endmodule