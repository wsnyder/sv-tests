/*
:name: fx68k
:description: Full fx68k core test
:files: /home/travis/build/SymbiFlow/sv-tests/third_party/cores/fx68k/fx68k.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/fx68k/fx68kAlu.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/fx68k/uaddrPla.sv 
:should_fail: 0
:tags: fx68k
*/
