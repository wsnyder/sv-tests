/*
:name: wait_order
:description: The 'wait_order' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit wait_order;
endmodule