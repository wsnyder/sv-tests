/*
:name: until_with
:description: The 'until_with' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit until_with;
endmodule