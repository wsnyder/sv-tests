/*
:name: integer_unsigned_shortint
:description: shortint unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
shortint unsigned v;
endmodule