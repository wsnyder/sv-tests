/*
:name: integer_signed_int
:description: int signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
int signed v;
endmodule