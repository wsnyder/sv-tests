/*
:name: net_wor
:description: wor net test
:should_fail: 0
:tags: 6.6.3
*/
module top();
wor v;
endmodule