/*
:name: net_supply1
:description: supply1 net test
:should_fail: 0
:tags: 6.6.6
*/
module top();
supply1 v;
endmodule