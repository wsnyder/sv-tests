/*
:name: net_supply0
:description: supply0 net test
:should_fail: 0
:tags: 6.6.6
*/
module top();
supply0 v;
endmodule