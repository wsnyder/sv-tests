/*
:name: s_until
:description: The 's_until' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit s_until;
endmodule