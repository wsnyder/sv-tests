/*
:name: supply0
:description: The 'supply0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit supply0;
endmodule