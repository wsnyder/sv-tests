/*
:name: pulsestyle_ondetect
:description: The 'pulsestyle_ondetect' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit pulsestyle_ondetect;
endmodule