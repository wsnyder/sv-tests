/*
:name: notif0
:description: The 'notif0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit notif0;
endmodule