/*
:name: always_latch
:description: The 'always_latch' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit always_latch;
endmodule