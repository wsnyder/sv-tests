/*
:name: net_triand
:description: triand net test
:should_fail: 0
:tags: 6.6.3
*/
module top();
triand v;
endmodule