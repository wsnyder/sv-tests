/*
:name: ibex
:description: Full ibex core test
:files: /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/examples/sim/rtl/prim_clock_gating.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_pkg.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_alu.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_compressed_decoder.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_controller.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_cs_registers.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_decoder.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_ex_block.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_id_stage.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_if_stage.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_load_store_unit.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_multdiv_slow.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_multdiv_fast.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_prefetch_buffer.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_fetch_fifo.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_pmp.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_core.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl/ibex_register_file_ff.sv 
:incdirs: /home/travis/build/SymbiFlow/sv-tests/third_party/cores/ibex/rtl 
:should_fail: 0
:tags: ibex
*/
