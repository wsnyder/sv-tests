/*
:name: endchecker
:description: The 'endchecker' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit endchecker;
endmodule