/*
:name: always_comb
:description: The 'always_comb' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit always_comb;
endmodule