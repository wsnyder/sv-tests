/*
:name: weak0
:description: The 'weak0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit weak0;
endmodule