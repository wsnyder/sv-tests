/*
:name: integer_bit
:description: bit net test
:should_fail: 0
:tags: 6.11
*/
module top();
bit v;
endmodule