/*
:name: join_any
:description: The 'join_any' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit join_any;
endmodule