/*
:name: integer_time
:description: time net test
:should_fail: 0
:tags: 6.11
*/
module top();
time v;
endmodule