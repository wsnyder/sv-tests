/*
:name: integer_unsigned_integer
:description: integer unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
integer unsigned v;
endmodule