/*
:name: swerv
:description: Full swerv core test
:files: /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/configs/snapshots/default/common_defines.vh /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/include/build.h /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/include/global.h /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/include/swerv_types.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/swerv_wrapper.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/mem.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/pic_ctrl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/swerv.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dma_ctrl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_aln_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_compress_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_ifc_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_bp_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_ic_mem.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_mem_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu_iccm_mem.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/ifu/ifu.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec_decode_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec_gpr_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec_ib_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec_tlu_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec_trigger.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dec/dec.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/exu/exu_alu_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/exu/exu_mul_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/exu/exu_div_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/exu/exu.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_clkdomain.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_addrcheck.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_lsc_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_stbuf.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_bus_buffer.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_bus_intf.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_ecc.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_dccm_mem.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_dccm_ctl.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lsu/lsu_trigger.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dbg/dbg.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dmi/dmi_wrapper.v /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dmi/dmi_jtag_to_core_sync.v /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dmi/rvjtag_tap.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lib/beh_lib.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lib/mem_lib.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lib/ahb_to_axi4.sv /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lib/axi4_to_ahb.sv 
:incdirs: /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/include /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/lib /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/design/dmi /home/travis/build/SymbiFlow/sv-tests/third_party/cores/swerv/configs/snapshots/default 
:should_fail: 0
:tags: swerv
:top_module: swerv_wrapper
*/
