/*
:name: s_always
:description: The 's_always' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit s_always;
endmodule