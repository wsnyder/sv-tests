/*
:name: integer_signed_longint
:description: longint signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
longint signed v;
endmodule