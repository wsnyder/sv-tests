/*
:name: shortreal
:description: The 'shortreal' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit shortreal;
endmodule