/*
:name: integer_byte
:description: byte net test
:should_fail: 0
:tags: 6.11
*/
module top();
byte v;
endmodule