/*
:name: notif1
:description: The 'notif1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit notif1;
endmodule