/*
:name: and_assignment
:description: &= assignment test
:should_fail: 0
:tags: 11.4.1
*/
module top();
int a = 12;
int b = 5;
initial begin
    a &= b;
end
endmodule