/*
:name: chandle
:description: The 'chandle' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit chandle;
endmodule