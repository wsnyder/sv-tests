/*
:name: highz0
:description: The 'highz0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit highz0;
endmodule