/*
:name: until
:description: The 'until' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit until;
endmodule