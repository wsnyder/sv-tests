/*
:name: supply1
:description: The 'supply1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit supply1;
endmodule