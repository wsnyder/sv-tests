/*
:name: s_nexttime
:description: The 's_nexttime' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit s_nexttime;
endmodule