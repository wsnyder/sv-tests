/*
:name: weak1
:description: The 'weak1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit weak1;
endmodule