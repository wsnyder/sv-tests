/*
:name: tri1
:description: The 'tri1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit tri1;
endmodule