/*
:name: integer_unsigned_byte
:description: byte unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
byte unsigned v;
endmodule