/*
:name: integer_logic
:description: logic net test
:should_fail: 0
:tags: 6.11
*/
module top();
logic v;
endmodule