/*
:name: integer_reg
:description: reg net test
:should_fail: 0
:tags: 6.11
*/
module top();
reg v;
endmodule