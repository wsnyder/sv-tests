/*
:name: net_tri1
:description: tri1 net test
:should_fail: 0
:tags: 6.6.5
*/
module top();
tri1 v;
endmodule