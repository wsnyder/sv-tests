/*
:name: unique0
:description: The 'unique0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit unique0;
endmodule