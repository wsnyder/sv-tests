/*
:name: integer_unsigned_int
:description: int unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
int unsigned v;
endmodule