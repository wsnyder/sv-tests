/*
:name: and
:description: The 'and' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit and;
endmodule