/*
:name: s_eventually
:description: The 's_eventually' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit s_eventually;
endmodule