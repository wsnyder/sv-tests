/*
:name: integer_unsigned_reg
:description: reg unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
reg unsigned v;
endmodule