/*
:name: s_until_with
:description: The 's_until_with' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit s_until_with;
endmodule