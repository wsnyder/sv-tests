/*
:name: highz1
:description: The 'highz1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit highz1;
endmodule