/*
:name: tri
:description: The 'tri' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit tri;
endmodule