/*
:name: strong1
:description: The 'strong1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit strong1;
endmodule