/*
:name: integer_unsigned_time
:description: time unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
time unsigned v;
endmodule