/*
:name: defparam
:description: The 'defparam' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit defparam;
endmodule