/*
:name: specify
:description: The 'specify' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit specify;
endmodule