/*
:name: integer_signed_reg
:description: reg signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
reg signed v;
endmodule