/*
:name: pull1
:description: The 'pull1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit pull1;
endmodule