/*
:name: integer_shortint
:description: shortint net test
:should_fail: 0
:tags: 6.11
*/
module top();
shortint v;
endmodule