/*
:name: net_trireg
:description: trireg net test
:should_fail: 0
:tags: 6.6.4
*/
module top();
trireg v;
endmodule