/*
:name: net_tri0
:description: tri0 net test
:should_fail: 0
:tags: 6.6.5
*/
module top();
tri0 v;
endmodule