/*
:name: integer_unsigned_logic
:description: logic unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
logic unsigned v;
endmodule