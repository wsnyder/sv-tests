/*
:name: sync_accept_on
:description: The 'sync_accept_on' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit sync_accept_on;
endmodule