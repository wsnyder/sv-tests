/*
:name: net_wire
:description: wire net test
:should_fail: 0
:tags: 6.6.1
*/
module top();
wire v;
endmodule