/*
:name: integer_unsigned_bit
:description: bit unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
bit unsigned v;
endmodule