/*
:name: tranif1
:description: The 'tranif1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit tranif1;
endmodule