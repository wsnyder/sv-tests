/*
:name: join_none
:description: The 'join_none' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit join_none;
endmodule