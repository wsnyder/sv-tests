/*
:name: bufif0
:description: The 'bufif0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit bufif0;
endmodule