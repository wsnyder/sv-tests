/*
:name: tranif0
:description: The 'tranif0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit tranif0;
endmodule