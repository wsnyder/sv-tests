/*
:name: ignore_bins
:description: The 'ignore_bins' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit ignore_bins;
endmodule