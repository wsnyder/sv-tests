/*
:name: net_uwire
:description: uwire net test
:should_fail: 0
:tags: 6.6.2
*/
module top();
uwire v;
endmodule