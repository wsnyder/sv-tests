/*
:name: rtranif1
:description: The 'rtranif1' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit rtranif1;
endmodule