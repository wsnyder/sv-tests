/*
:name: reject_on
:description: The 'reject_on' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit reject_on;
endmodule