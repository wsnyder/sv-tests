/*
:name: tri0
:description: The 'tri0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit tri0;
endmodule