/*
:name: integer_signed_logic
:description: logic signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
logic signed v;
endmodule