/*
:name: integer_signed_shortint
:description: shortint signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
shortint signed v;
endmodule