/*
:name: sync_reject_on
:description: The 'sync_reject_on' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit sync_reject_on;
endmodule