/*
:name: always_ff
:description: The 'always_ff' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit always_ff;
endmodule