/*
:name: output
:description: The 'output' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit output;
endmodule