/*
:name: strong0
:description: The 'strong0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit strong0;
endmodule