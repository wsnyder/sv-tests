/*
:name: global
:description: The 'global' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit global;
endmodule