/*
:name: net_trior
:description: trior net test
:should_fail: 0
:tags: 6.6.3
*/
module top();
trior v;
endmodule