/*
:name: rtran
:description: The 'rtran' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit rtran;
endmodule