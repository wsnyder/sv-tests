/*
:name: net_tri
:description: tri net test
:should_fail: 0
:tags: 6.6.1
*/
module top();
tri v;
endmodule