/*
:name: integer_int
:description: int net test
:should_fail: 0
:tags: 6.11
*/
module top();
int v;
endmodule