/*
:name: integer_unsigned_longint
:description: longint unsigned net test
:should_fail: 0
:tags: 6.11
*/
module top();
longint unsigned v;
endmodule