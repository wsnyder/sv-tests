/*
:name: integer_signed_integer
:description: integer signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
integer signed v;
endmodule