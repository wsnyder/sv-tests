/*
:name: intersect
:description: The 'intersect' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit intersect;
endmodule