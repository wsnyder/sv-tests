/*
:name: integer_longint
:description: longint net test
:should_fail: 0
:tags: 6.11
*/
module top();
longint v;
endmodule