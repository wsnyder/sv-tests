/*
:name: rtranif0
:description: The 'rtranif0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit rtranif0;
endmodule