/*
:name: nor
:description: The 'nor' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit nor;
endmodule