/*
:name: integer_signed_time
:description: time signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
time signed v;
endmodule