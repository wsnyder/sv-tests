/*
:name: integer_integer
:description: integer net test
:should_fail: 0
:tags: 6.11
*/
module top();
integer v;
endmodule