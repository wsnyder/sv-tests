/*
:name: illegal_bins
:description: The 'illegal_bins' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit illegal_bins;
endmodule