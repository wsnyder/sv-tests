/*
:name: accept_on
:description: The 'accept_on' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit accept_on;
endmodule