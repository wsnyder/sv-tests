/*
:name: endprogram
:description: The 'endprogram' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit endprogram;
endmodule