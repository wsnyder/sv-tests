/*
:name: integer_signed_byte
:description: byte signed net test
:should_fail: 0
:tags: 6.11
*/
module top();
byte signed v;
endmodule