/*
:name: endcase
:description: The 'endcase' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit endcase;
endmodule