/*
:name: pull0
:description: The 'pull0' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit pull0;
endmodule