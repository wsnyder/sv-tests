/*
:name: time
:description: The 'time' keyword should be reserved
:should_fail: 1
:tags: 5.6.2
*/
module top();
    bit time;
endmodule